
`ifndef PredictionSignals
`define PredictionSignals



`define NOBRANCH            3'b000


`define NOGUESS_INCORRECT   3'b100
`define NOGUESS_CORRECT     3'b101

`define GUESS_INCORRECT     3'b110
`define GUESS_CORRECT       3'b111

`endif //OPCODE