/*
List of Register Names.
*/

`ifndef RegNames
`define ALUOP

`define x0  5'b00000
`define x1  5'b00001
`define x2  5'b00010
`define x3  5'b00011
`define x4  5'b00100
`define x5  5'b00101
`define x6  5'b00110
`define x7  5'b00111
`define x8  5'b01000
`define x9  5'b01001
`define x10 5'b01010
`define x11 5'b01011
`define x12 5'b01100
`define x13 5'b01101
`define x14 5'b01110
`define x15 5'b01111
`define x16 5'b10000
`define x17 5'b10001
`define x18 5'b10010
`define x19 5'b10011
`define x20 5'b10100
`define x21 5'b10101
`define x22 5'b10110
`define x23 5'b10111
`define x24 5'b11000
`define x25 5'b11001
`define x26 5'b11010
`define x27 5'b11011
`define x28 5'b11100
`define x29 5'b11101
`define x30 5'b11110
`define x31 5'b11111


`endif //RegNames
