/*
Module:
    Immediate Selector (ImmSel)

Description:
    This module is not necessasrily needed, since the instruction 
    is sent to the immediate generator to figure it out and can 
    be determined by that module.

Authors:
    Matthew Dharmawan and Reuben Koshy Thomas

*/